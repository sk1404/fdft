`timescale 1ns/1ps

module scan_dff_mux (
    input  wire D,     // Normal data input
    input  wire SD,    // Scan data input
    input  wire SE,    // Scan enable (mux select)
    input  wire CLK,   // Clock
    input  wire RST,   // Asynchronous active-high reset
    output reg  Q      // Output
);

    wire mux_out;

    // 2:1 MUX: If SE == 1, select SD; else select D
    assign mux_out = SE ? SD : D;

    // Positive-edge triggered DFF with async reset
    always @(posedge CLK or posedge RST) begin
        if (RST)
            Q <= 1'b0;
        else
            Q <= mux_out;
    end

endmodule


// Generated by Cadence Genus(TM) Synthesis Solution 20.10-p001_1
// Generated on: Jul 12 2025 15:27:44 IST (Jul 12 2025 09:57:44 UTC)

// Verification Directory fv/counter_4bit 

module counter_4bit(clk, reset, count,SD,SE);
  input clk, reset,SD,SE;
  output [3:0] count;
  wire clk, reset;
  wire [3:0] count;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8;

  //DFFHQX1 \count_reg[3] (.CK (clk), .D (n_8), .Q (count[3]));
  scan_dff_mux s4(.D(n_8),.SD(count[2]),.SE(SE),.CLK(clk),.RST(reset),.Q(count[3]));
  NOR2XL g60(.A (reset), .B (n_7), .Y (n_8));

  //DFFHQX1 \count_reg[2] (.CK (clk), .D (n_6), .Q (count[2]));
  scan_dff_mux s3(.D(n_6),.SD(count[1]),.SE(SE),.CLK(clk),.RST(reset),.Q(count[2])); 
 //DFFHQX1 \count_reg[1] (.CK (clk), .D (n_4), .Q (count[1]));
  scan_dff_mux s2(.D(n_4),.SD(count[0]),.SE(SE),.CLK(clk),.RST(reset),.Q(count[1]));
  XNOR2X1 g62(.A (n_5), .B (count[3]), .Y (n_7));
  AOI211XL g63(.A0 (n_1), .A1 (n_2), .B0 (reset), .C0 (n_5), .Y (n_6));
  NOR2XL g66(.A (reset), .B (n_3), .Y (n_4));
  OAI21XL g68(.A0 (count[0]), .A1 (count[1]), .B0 (n_2), .Y (n_3));
  NOR2XL g65(.A (n_1), .B (n_2), .Y (n_5));
  
  //DFFHQX1 \count_reg[0] (.CK (clk), .D (n_0), .Q (count[0]));
  scan_dff_mux s1(.D(n_0),.SD(SD),.SE(SE),.CLK(clk),.RST(reset),.Q(count[0]));
  NOR2XL g69(.A (reset), .B (count[0]), .Y (n_0));
  NAND2XL g70(.A (count[1]), .B (count[0]), .Y (n_2));
  INVXL g71(.A (count[2]), .Y (n_1));
endmodule


module counter_4bit_tb;

  // Inputs
  reg clk;
  reg reset;
  reg SD;
  reg SE;

  // Outputs
  wire [3:0] count;

  // Instantiate the Unit Under Test (UUT)
  counter_4bit uut (
    .clk(clk),
    .reset(reset),
    .count(count),
    .SD(SD),
    .SE(SE)
  );

  // Clock Generation: 10ns period
  initial clk = 0;
  always #5 clk = ~clk;

  // Test Sequence
  initial begin
    $display("Starting Testbench...");
    $dumpfile("counter_4bit.vcd");
    $dumpvars(0, counter_4bit_tb);

    // Initialize inputs
    reset = 1;
    SD = 0;
    SE = 0;

    // Apply reset
    #10;
    reset = 0;

    // Count normally (SE = 0)
    $display("Normal Counting...");
    repeat (16) begin
      #10;
      $display("Time = %0t | Count = %b", $time, count);
    end

    // Apply reset again
    reset = 1; #10;
    reset = 0; #10;

    // Scan mode operation
    SE = 1; // Enable scan mode
    $display("Scan Mode Operation...");
    SD = 1;
    #10;
    $display("Time = %0t | Count = %b (Scan Mode)", $time, count);
    
    SD = 0;
    #10;
    $display("Time = %0t | Count = %b (Scan Mode)", $time, count);

    SE = 0; // Return to normal mode

    // Final few clocks in normal mode
    $display("Return to Normal Counting...");
    repeat (5) begin
      #10;
      $display("Time = %0t | Count = %b", $time, count);
    end

    $finish;
  end

endmodule
